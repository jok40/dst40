/******************************************************************************

  Функция Fe для ядра DST40.

  Реализована полностью комбинаторно. Изначально было пять входов, но потом
  сократили до четырёх - выкинули младший вход, так как в исходной таблице
  все биты повторялись по два раза.

******************************************************************************/

module Fe
(
  input   [3:0] in,
  output        out
);

reg     i;
assign  out = i;

always  @( in )
begin
  case( in )
    4'b 0000: i = 0;
    4'b 0001: i = 1;
    4'b 0010: i = 0;
    4'b 0011: i = 1;
    4'b 0100: i = 0;
    4'b 0101: i = 0;
    4'b 0110: i = 1;
    4'b 0111: i = 1;
    4'b 1000: i = 1;
    4'b 1001: i = 1;
    4'b 1010: i = 0;
    4'b 1011: i = 0;
    4'b 1100: i = 1;
    4'b 1101: i = 0;
    4'b 1110: i = 1;
    default : i = 0;
  endcase
end

endmodule
