/******************************************************************************

  Функция Fc для ядра DST40.

  Реализована полностью комбинаторно.

******************************************************************************/

module Fc
(
  input   [4:0] in,
  output        out
);


reg     i;
assign  out = i;

always  @( in )
begin
  case( in )
    5'b 00000: i = 0;
    5'b 00001: i = 0;
    5'b 00010: i = 1;
    5'b 00011: i = 0;
    5'b 00100: i = 1;
    5'b 00101: i = 1;
    5'b 00110: i = 1;
    5'b 00111: i = 0;
    5'b 01000: i = 1;
    5'b 01001: i = 0;
    5'b 01010: i = 1;
    5'b 01011: i = 1;
    5'b 01100: i = 1;
    5'b 01101: i = 0;
    5'b 01110: i = 0;
    5'b 01111: i = 0;
    5'b 10000: i = 0;
    5'b 10001: i = 0;
    5'b 10010: i = 1;
    5'b 10011: i = 1;
    5'b 10100: i = 1;
    5'b 10101: i = 1;
    5'b 10110: i = 0;
    5'b 10111: i = 0;
    5'b 11000: i = 0;
    5'b 11001: i = 1;
    5'b 11010: i = 0;
    5'b 11011: i = 1;
    5'b 11100: i = 0;
    5'b 11101: i = 1;
    5'b 11110: i = 0;
    default  : i = 1;
  endcase
end

endmodule
