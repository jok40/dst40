/******************************************************************************

  Функция Fh для ядра DST40.

  Реализована полностью комбинаторно.

******************************************************************************/

module Fh
(
  input   [3:0] in,
  output  [1:0] out
);


reg [1:0] i;

assign  out = i;

always  @( in )
begin
  case( in )
    4'b 0000: i = 2'b 00;
    4'b 0001: i = 2'b 00;
    4'b 0010: i = 2'b 10;
    4'b 0011: i = 2'b 11;
    4'b 0100: i = 2'b 11;
    4'b 0101: i = 2'b 01;
    4'b 0110: i = 2'b 10;
    4'b 0111: i = 2'b 01;
    4'b 1000: i = 2'b 01;
    4'b 1001: i = 2'b 10;
    4'b 1010: i = 2'b 01;
    4'b 1011: i = 2'b 11;
    4'b 1100: i = 2'b 11;
    4'b 1101: i = 2'b 10;
    4'b 1110: i = 2'b 00;
    default : i = 2'b 00;
  endcase
end


endmodule
